module fifo_integrity();
endmodule